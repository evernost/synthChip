-- ============================================================================
-- Project        : synthChip
-- Module name    : synthChip_pkg
-- File name      : synthChip_pkg.vhd
-- File type      : VHDL 2008
-- Purpose        : package definition for the synthChip FPGA
-- Author         : QuBi (nitrogenium@outlook.fr)
-- Creation date  : August 6th, 2025
-- ----------------------------------------------------------------------------
-- Best viewed with space indentation (2 spaces)
-- ============================================================================

-- ============================================================================
-- CONTENT IS GENERATED AUTOMATICALLY USING 'makeFPGA.tcl'
-- ! DO NOT MODIFY IT !
-- ============================================================================

-- ============================================================================
-- LIBRARIES
-- ============================================================================
-- Standard libraries
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;



-- ============================================================================
-- PACKAGE DESCRIPTION
-- ============================================================================
package synthChip_pkg is
  
  -- --------------------------------------------------------------------------
  -- Constants / Types
  -- --------------------------------------------------------------------------
  constant FPGA_VERSION  : STD_LOGIC_VECTOR(31 downto 0) := 1;
  
  
  -- --------------------------------------------------------------------------
  -- Components
  -- --------------------------------------------------------------------------
  -- None.
  
end package synthChip_pkg;
  
  
  
-- ============================================================================
-- PACKAGE DESCRIPTION
-- ============================================================================
package body synthChip_pkg is 
  
  -- None.
  
end package body;
