-- ============================================================================
-- Project        : Blinky
-- Module name    : blinky
-- File name      : blinky.vhd
-- File type      : VHDL 2008
-- Purpose        : package definition for the Blinky module
-- Author         : QuBi (nitrogenium@outlook.fr)
-- Creation date  : August 11, 2025 at 00:14
-- ----------------------------------------------------------------------------
-- Best viewed with space indentation (2 spaces)
-- ============================================================================

-- ============================================================================
-- CONTENT IS GENERATED AUTOMATICALLY USING 'makeBrightnessLut.py'.
-- ! DO NOT MODIFY IT !
-- ============================================================================

-- ============================================================================
-- LIBRARIES
-- ============================================================================
-- Standard libraries
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;



-- ============================================================================
-- PACKAGE DESCRIPTION
-- ============================================================================
package blinky_pkg is
  
  -- --------------------------------------------------------------------------
  -- Constants / Types
  -- --------------------------------------------------------------------------
  constant PWM_RESOL_NBITS  : INTEGER := 9;
  constant BRIGHTNESS_STEPS : INTEGER := 128;
  
  type ROM_TYPE is array (0 to (BRIGHTNESS_STEPS-1)) of STD_LOGIC_VECTOR((PWM_RESOL_NBITS-1) downto 0);
 
  constant BRIGHTNESS_ROM : ROM_TYPE := 
  (
    0 => "000000000",    -- PWM(0) = 0/512
    1 => "000000000",    -- PWM(1) = 0/512
    2 => "000000000",    -- PWM(2) = 0/512
    3 => "000000000",    -- PWM(3) = 0/512
    4 => "000000000",    -- PWM(4) = 0/512
    5 => "000000000",    -- PWM(5) = 0/512
    6 => "000000000",    -- PWM(6) = 0/512
    7 => "000000000",    -- PWM(7) = 0/512
    8 => "000000000",    -- PWM(8) = 0/512
    9 => "000000001",    -- PWM(9) = 1/512
    10 => "000000001",    -- PWM(10) = 1/512
    11 => "000000001",    -- PWM(11) = 1/512
    12 => "000000001",    -- PWM(12) = 1/512
    13 => "000000001",    -- PWM(13) = 1/512
    14 => "000000001",    -- PWM(14) = 1/512
    15 => "000000001",    -- PWM(15) = 1/512
    16 => "000000001",    -- PWM(16) = 1/512
    17 => "000000001",    -- PWM(17) = 1/512
    18 => "000000001",    -- PWM(18) = 1/512
    19 => "000000010",    -- PWM(19) = 2/512
    20 => "000000010",    -- PWM(20) = 2/512
    21 => "000000010",    -- PWM(21) = 2/512
    22 => "000000010",    -- PWM(22) = 2/512
    23 => "000000010",    -- PWM(23) = 2/512
    24 => "000000010",    -- PWM(24) = 2/512
    25 => "000000010",    -- PWM(25) = 2/512
    26 => "000000011",    -- PWM(26) = 3/512
    27 => "000000011",    -- PWM(27) = 3/512
    28 => "000000011",    -- PWM(28) = 3/512
    29 => "000000011",    -- PWM(29) = 3/512
    30 => "000000011",    -- PWM(30) = 3/512
    31 => "000000100",    -- PWM(31) = 4/512
    32 => "000000100",    -- PWM(32) = 4/512
    33 => "000000100",    -- PWM(33) = 4/512
    34 => "000000100",    -- PWM(34) = 4/512
    35 => "000000101",    -- PWM(35) = 5/512
    36 => "000000101",    -- PWM(36) = 5/512
    37 => "000000101",    -- PWM(37) = 5/512
    38 => "000000101",    -- PWM(38) = 5/512
    39 => "000000110",    -- PWM(39) = 6/512
    40 => "000000110",    -- PWM(40) = 6/512
    41 => "000000110",    -- PWM(41) = 6/512
    42 => "000000111",    -- PWM(42) = 7/512
    43 => "000000111",    -- PWM(43) = 7/512
    44 => "000001000",    -- PWM(44) = 8/512
    45 => "000001000",    -- PWM(45) = 8/512
    46 => "000001000",    -- PWM(46) = 8/512
    47 => "000001001",    -- PWM(47) = 9/512
    48 => "000001001",    -- PWM(48) = 9/512
    49 => "000001010",    -- PWM(49) = 10/512
    50 => "000001010",    -- PWM(50) = 10/512
    51 => "000001011",    -- PWM(51) = 11/512
    52 => "000001100",    -- PWM(52) = 12/512
    53 => "000001100",    -- PWM(53) = 12/512
    54 => "000001101",    -- PWM(54) = 13/512
    55 => "000001110",    -- PWM(55) = 14/512
    56 => "000001110",    -- PWM(56) = 14/512
    57 => "000001111",    -- PWM(57) = 15/512
    58 => "000010000",    -- PWM(58) = 16/512
    59 => "000010001",    -- PWM(59) = 17/512
    60 => "000010010",    -- PWM(60) = 18/512
    61 => "000010011",    -- PWM(61) = 19/512
    62 => "000010100",    -- PWM(62) = 20/512
    63 => "000010101",    -- PWM(63) = 21/512
    64 => "000010110",    -- PWM(64) = 22/512
    65 => "000010111",    -- PWM(65) = 23/512
    66 => "000011000",    -- PWM(66) = 24/512
    67 => "000011001",    -- PWM(67) = 25/512
    68 => "000011010",    -- PWM(68) = 26/512
    69 => "000011100",    -- PWM(69) = 28/512
    70 => "000011101",    -- PWM(70) = 29/512
    71 => "000011111",    -- PWM(71) = 31/512
    72 => "000100000",    -- PWM(72) = 32/512
    73 => "000100010",    -- PWM(73) = 34/512
    74 => "000100100",    -- PWM(74) = 36/512
    75 => "000100110",    -- PWM(75) = 38/512
    76 => "000101000",    -- PWM(76) = 40/512
    77 => "000101010",    -- PWM(77) = 42/512
    78 => "000101100",    -- PWM(78) = 44/512
    79 => "000101110",    -- PWM(79) = 46/512
    80 => "000110000",    -- PWM(80) = 48/512
    81 => "000110011",    -- PWM(81) = 51/512
    82 => "000110101",    -- PWM(82) = 53/512
    83 => "000111000",    -- PWM(83) = 56/512
    84 => "000111011",    -- PWM(84) = 59/512
    85 => "000111110",    -- PWM(85) = 62/512
    86 => "001000001",    -- PWM(86) = 65/512
    87 => "001000100",    -- PWM(87) = 68/512
    88 => "001001000",    -- PWM(88) = 72/512
    89 => "001001100",    -- PWM(89) = 76/512
    90 => "001001111",    -- PWM(90) = 79/512
    91 => "001010011",    -- PWM(91) = 83/512
    92 => "001011000",    -- PWM(92) = 88/512
    93 => "001011100",    -- PWM(93) = 92/512
    94 => "001100001",    -- PWM(94) = 97/512
    95 => "001100110",    -- PWM(95) = 102/512
    96 => "001101011",    -- PWM(96) = 107/512
    97 => "001110000",    -- PWM(97) = 112/512
    98 => "001110110",    -- PWM(98) = 118/512
    99 => "001111100",    -- PWM(99) = 124/512
    100 => "010000010",    -- PWM(100) = 130/512
    101 => "010001000",    -- PWM(101) = 136/512
    102 => "010001111",    -- PWM(102) = 143/512
    103 => "010010110",    -- PWM(103) = 150/512
    104 => "010011110",    -- PWM(104) = 158/512
    105 => "010100110",    -- PWM(105) = 166/512
    106 => "010101110",    -- PWM(106) = 174/512
    107 => "010110111",    -- PWM(107) = 183/512
    108 => "011000000",    -- PWM(108) = 192/512
    109 => "011001010",    -- PWM(109) = 202/512
    110 => "011010100",    -- PWM(110) = 212/512
    111 => "011011111",    -- PWM(111) = 223/512
    112 => "011101010",    -- PWM(112) = 234/512
    113 => "011110101",    -- PWM(113) = 245/512
    114 => "100000010",    -- PWM(114) = 258/512
    115 => "100001111",    -- PWM(115) = 271/512
    116 => "100011100",    -- PWM(116) = 284/512
    117 => "100101011",    -- PWM(117) = 299/512
    118 => "100111001",    -- PWM(118) = 313/512
    119 => "101001001",    -- PWM(119) = 329/512
    120 => "101011010",    -- PWM(120) = 346/512
    121 => "101101011",    -- PWM(121) = 363/512
    122 => "101111101",    -- PWM(122) = 381/512
    123 => "110010000",    -- PWM(123) = 400/512
    124 => "110100100",    -- PWM(124) = 420/512
    125 => "110111001",    -- PWM(125) = 441/512
    126 => "111001111",    -- PWM(126) = 463/512
    127 => "111100111"     -- PWM(127) = 487/512
  );
  
  -- --------------------------------------------------------------------------
  -- Components
  -- --------------------------------------------------------------------------
  -- None.
  
end package blinky_pkg;
  
  
  
-- ============================================================================
-- PACKAGE DESCRIPTION
-- ============================================================================
package body blinky_pkg is 
  
  -- None.
  
end package body;
